// turn off that dm led
// Author: Mikhail w/ the help of Ryan 
// 2/1/2025
//////////////////////////////////////////////////////////////////////////

module whiteOut (
   output logic red, green, blue
);
   assign red = 0;
   assign blue = 0;
   assign green = 0;
endmodule
